library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mux is
    Port ( SEL : in  STD_LOGIC;
           IN1  : in  STD_LOGIC;
           IN2   : in  STD_LOGIC;
           outM   : out STD_LOGIC);
end mux;

architecture Behavioral of mux is
begin
    outM <=  IN1 when (SEL = '0') else IN2;
end Behavioral;
